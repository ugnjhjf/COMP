
module And_Or_Latch(
    input set,reset,
    output data)

assign 


endmodule